

module enRoundKey(dataa, datab, result);
  input [31:0] dataa, datab;
  output [31:0] result;



endmodule
